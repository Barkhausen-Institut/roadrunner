localparam WORLD = "Welt";