localparam HELLO = "Hallo";