module m1;

endmodule