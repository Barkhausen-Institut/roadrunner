////    ////////////
////    ////////////
////
////
////////////    ////
////////////    ////
////    ////    ////
////    ////    ////
////////////
////////////


module SimTest();

import "DPI-C" function void DPIGreeting();
import "DPI-C" function void DPISuccess();
import RREnv::*;

initial DPIGreeting();

initial DPISuccess();

endmodule