module mod2;

endmodule